module xillybus_core
  (
  input  M_AXI_ACP_ARREADY_w,
  input  M_AXI_ACP_AWREADY_w,
  input [1:0] M_AXI_ACP_BRESP_w,
  input  M_AXI_ACP_BVALID_w,
  input [63:0] M_AXI_ACP_RDATA_w,
  input  M_AXI_ACP_RLAST_w,
  input [1:0] M_AXI_ACP_RRESP_w,
  input  M_AXI_ACP_RVALID_w,
  input  M_AXI_ACP_WREADY_w,
  input [31:0] S_AXI_ARADDR_w,
  input  S_AXI_ARVALID_w,
  input [31:0] S_AXI_AWADDR_w,
  input  S_AXI_AWVALID_w,
  input  S_AXI_BREADY_w,
  input  S_AXI_RREADY_w,
  input [31:0] S_AXI_WDATA_w,
  input [3:0] S_AXI_WSTRB_w,
  input  S_AXI_WVALID_w,
  input  bus_clk_w,
  input  bus_rst_n_w,
  input [31:0] user_r_accx_read_data_w,
  input  user_r_accx_read_empty_w,
  input  user_r_accx_read_eof_w,
  input [31:0] user_r_accy_read_data_w,
  input  user_r_accy_read_empty_w,
  input  user_r_accy_read_eof_w,
  input [31:0] user_r_accz_read_data_w,
  input  user_r_accz_read_empty_w,
  input  user_r_accz_read_eof_w,
  input [31:0] user_r_gyrox_read_data_w,
  input  user_r_gyrox_read_empty_w,
  input  user_r_gyrox_read_eof_w,
  input [31:0] user_r_gyroy_read_data_w,
  input  user_r_gyroy_read_empty_w,
  input  user_r_gyroy_read_eof_w,
  input [31:0] user_r_gyroz_read_data_w,
  input  user_r_gyroz_read_empty_w,
  input  user_r_gyroz_read_eof_w,
  input [31:0] user_r_magx_read_data_w,
  input  user_r_magx_read_empty_w,
  input  user_r_magx_read_eof_w,
  input [31:0] user_r_magy_read_data_w,
  input  user_r_magy_read_empty_w,
  input  user_r_magy_read_eof_w,
  input [31:0] user_r_magz_read_data_w,
  input  user_r_magz_read_empty_w,
  input  user_r_magz_read_eof_w,
  input [31:0] user_r_op_data_w,
  input  user_r_op_empty_w,
  input  user_r_op_eof_w,
  input [31:0] user_r_qa_read_data_w,
  input  user_r_qa_read_empty_w,
  input  user_r_qa_read_eof_w,
  input [31:0] user_r_qb_read_data_w,
  input  user_r_qb_read_empty_w,
  input  user_r_qb_read_eof_w,
  input [31:0] user_r_qc_read_data_w,
  input  user_r_qc_read_empty_w,
  input  user_r_qc_read_eof_w,
  input [31:0] user_r_qs_read_data_w,
  input  user_r_qs_read_empty_w,
  input  user_r_qs_read_eof_w,
  input  user_w_op_full_w,
  output [3:0] GPIO_LED_w,
  output [31:0] M_AXI_ACP_ARADDR_w,
  output [1:0] M_AXI_ACP_ARBURST_w,
  output [3:0] M_AXI_ACP_ARCACHE_w,
  output [3:0] M_AXI_ACP_ARLEN_w,
  output [2:0] M_AXI_ACP_ARPROT_w,
  output [2:0] M_AXI_ACP_ARSIZE_w,
  output  M_AXI_ACP_ARVALID_w,
  output [31:0] M_AXI_ACP_AWADDR_w,
  output [1:0] M_AXI_ACP_AWBURST_w,
  output [3:0] M_AXI_ACP_AWCACHE_w,
  output [3:0] M_AXI_ACP_AWLEN_w,
  output [2:0] M_AXI_ACP_AWPROT_w,
  output [2:0] M_AXI_ACP_AWSIZE_w,
  output  M_AXI_ACP_AWVALID_w,
  output  M_AXI_ACP_BREADY_w,
  output  M_AXI_ACP_RREADY_w,
  output [63:0] M_AXI_ACP_WDATA_w,
  output  M_AXI_ACP_WLAST_w,
  output [7:0] M_AXI_ACP_WSTRB_w,
  output  M_AXI_ACP_WVALID_w,
  output  S_AXI_ARREADY_w,
  output  S_AXI_AWREADY_w,
  output [1:0] S_AXI_BRESP_w,
  output  S_AXI_BVALID_w,
  output [31:0] S_AXI_RDATA_w,
  output [1:0] S_AXI_RRESP_w,
  output  S_AXI_RVALID_w,
  output  S_AXI_WREADY_w,
  output  host_interrupt_w,
  output  quiesce_w,
  output  user_r_accx_read_open_w,
  output  user_r_accx_read_rden_w,
  output  user_r_accy_read_open_w,
  output  user_r_accy_read_rden_w,
  output  user_r_accz_read_open_w,
  output  user_r_accz_read_rden_w,
  output  user_r_gyrox_read_open_w,
  output  user_r_gyrox_read_rden_w,
  output  user_r_gyroy_read_open_w,
  output  user_r_gyroy_read_rden_w,
  output  user_r_gyroz_read_open_w,
  output  user_r_gyroz_read_rden_w,
  output  user_r_magx_read_open_w,
  output  user_r_magx_read_rden_w,
  output  user_r_magy_read_open_w,
  output  user_r_magy_read_rden_w,
  output  user_r_magz_read_open_w,
  output  user_r_magz_read_rden_w,
  output  user_r_op_open_w,
  output  user_r_op_rden_w,
  output  user_r_qa_read_open_w,
  output  user_r_qa_read_rden_w,
  output  user_r_qb_read_open_w,
  output  user_r_qb_read_rden_w,
  output  user_r_qc_read_open_w,
  output  user_r_qc_read_rden_w,
  output  user_r_qs_read_open_w,
  output  user_r_qs_read_rden_w,
  output [31:0] user_w_op_data_w,
  output  user_w_op_open_w,
  output  user_w_op_wren_w
);
endmodule
